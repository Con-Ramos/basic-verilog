module mux_always #(parameter integer WIDTH = 1)(  //modulo mux realiza a selecao dos dados
    input wire [WIDTH-1:0] in_A,            //entrada 0, in_A = primeira entrada do mux
    input wire [WIDTH-1:0] in_B,            //entrada 1, in_B = segunda entrada do mux
    input wire sel,                         //sinal de selecao, qual das duas entradas sera passada para a saida
    output reg[WIDTH-1:0] mux_output  );    //saida do mux

    always @(*) //executa sempre que qualquer uma das entradas de um bloco combinacional ou sequencial muda de valor
        begin
            if (sel == 1)                   //se sel for 1(true) a saida sera igual a in_B
                mux_output = in_B;
            else                            //se nao, (false) a saida sera igual a in_A
                mux_output = in_A;
        end
endmodule                                   //final do modulo
